D:\Proyectos\Texturas\TxEstudio 2.0 (Enero2010)\TxEstudioApplication\bin\Debug\
7.bmp
D:\Proyectos\Texturas\TxEstudio 2.0 (Enero2010)\TxEstudioApplication\bin\Debug\
10.bmp
D:\Proyectos\Texturas\TxEstudio 2.0 (Enero2010)\TxEstudioApplication\bin\Debug\
som.bmp
D:\Proyectos\Texturas\TxEstudio 2.0 (Enero2010)\TxEstudioApplication\bin\Debug\
Leopard1..bmp
D:\Proyectos\Texturas\TxEstudio 2.0 (Enero2010)\TxEstudioApplication\bin\Debug\
0.jpg
D:\Proyectos\Proyecto TxEstudio\Union\TxEstudio 2.0 (Octubre)\TxEstudioApplication\bin\Debug\
2.bmp
D:\Buzon\Images\
mosaic_01_gt.bmp
D:\Buzon\Images\
mosaic_01_test.bmp
D:\Buzon\TxEstudio 2.0 (diciembre)\TxEstudioApplication\bin\Debug\
0.bmp
p
ebug\
0.bmp
lication\bin\Debug\
3.bmp
D:\ImagenesPrueba\Grafos\
E.bmp
ados Obtenidos\11 Plataforma TxEstudio Vers2\DemoTx\01 SegmRegiones\SWA\
Leon-SWA-Historia.bmp
btenidos\12 Bordes de Textura\5T\
5T+ts_mhs(5,15).bmp
sultados Obtenidos\12 Bordes de Textura\5T\
5T+gab_energ(4,22.5).bmp
nidos\12 Bordes de Textura\5T\
5T+gab_energ(4,0).bmp
D:\JLGil\Proyecto 2006\Proy. Segmentacion de Textura\Resultados Obtenidos\12 Bordes de Textura\5T\
5T+fo_min(7,7).bmp
